library ieee;
use ieee.std_logic_1164.all;

entity Test1top is
port (
    led : out std_logic_vector(15 downto 0)
);
end Test1top;

architecture rtl of Test1top is
begin
    led <= "0111111111010001";
end rtl;