library IEEE;
use ieee.std_logic_1164.all;

entity AND2_gate is
 port (
  X0, X1 : in std_logic;
  O : out std_logic
  ); 
end AND2_gate;

architecture rtl of AND2_gate is
begin
 O <= X1 and X0;
end rtl;